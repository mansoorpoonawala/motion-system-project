library ieee;
use ieee.std_logic_1164.all;

entity top_module is
    port (
        -- Clock and Reset
        sys_clk      : in  std_logic; -- 125MHz system clock from Zybo Z7
        sys_reset    : in  std_logic; -- System reset input (e.g., from a button)

        -- SPI Interface to ADXL345 (Connect to Pmod pins)
        spi_sclk_pin : out std_logic; -- SPI Serial Clock output
        spi_mosi_pin : out std_logic; -- SPI Master Out Slave In output
        spi_miso_pin : in  std_logic; -- SPI Master In Slave Out input
        spi_cs_pin   : out std_logic; -- SPI Chip Select output

        -- User LEDs on Zybo Z7
        leds         : out std_logic_vector(3 downto 0) -- Output to the 4 user LEDs
    );
end entity top_module;

architecture structural of top_module is

    -- Internal signals to connect modules
    signal clk_4mhz     : std_logic; -- 4MHz clock generated by iclk_gen
    signal acl_data_int : std_logic_vector(47 downto 0); -- Accelerometer data from spi_master (X, Y, Z - 16 bits each)
    signal spi_busy_int : std_logic; -- Signal indicating if SPI master is busy

    -- Component declarations for the modules to be instantiated
    -- These declarations must match the entity ports of the respective modules

    component iclk_gen
        port (
            clk       : in  std_logic; -- 125MHz input clock
            clk_4MHz  : out std_logic  -- 4MHz output clock
        );
    end component;

    component spi_master
        port (
            iclk       : in  std_logic; -- 4MHz clock input
            reset      : in  std_logic; -- Synchronous reset input
            miso       : in  std_logic; -- SPI Master In Slave Out
            sclk       : out std_logic; -- SPI Serial Clock (1MHz generated internally)
            mosi       : out std_logic; -- SPI Master Out Slave In
            cs         : out std_logic; -- SPI Chip Select (active low)
            acl_data   : out std_logic_vector(47 downto 0); -- Output accelerometer data (X[15:0], Y[15:0], Z[15:0])
            spi_busy   : out std_logic -- Indicates if SPI is busy
        );
    end component;

    component acl_led_indicator
        port (
            clk_125mhz : in  std_logic; -- 125MHz system clock
            reset      : in  std_logic; -- Synchronous reset input
            acl_data   : in  std_logic_vector(47 downto 0); -- Input accelerometer data

            leds_out   : out std_logic_vector(3 downto 0) -- Output to the 4 user LEDs
        );
    end component;

begin

    -- Instantiate the 4MHz clock generator
    iclk_gen_inst : iclk_gen
        port map (
            clk      => sys_clk,      -- Connect to the 125MHz system clock
            clk_4MHz => clk_4mhz      -- Connect to the internal 4MHz signal
        );

    -- Instantiate the SPI Master module
    spi_master_inst : spi_master
        port map (
            iclk       => clk_4mhz,     -- Connect to the generated 4MHz clock
            reset      => sys_reset,    -- Connect to the system reset
            miso       => spi_miso_pin, -- Connect to the physical MISO pin
            sclk       => spi_sclk_pin, -- Connect to the physical SCLK pin
            mosi       => spi_mosi_pin, -- Connect to the physical MOSI pin
            cs         => spi_cs_pin,   -- Connect to the physical CS pin
            acl_data   => acl_data_int, -- Connect to the internal accelerometer data signal
            spi_busy   => spi_busy_int  -- Connect to the internal SPI busy signal
        );

    -- Instantiate the Accelerometer Data LED Indicator module
    acl_led_indicator_inst : acl_led_indicator
        port map (
            clk_125mhz => sys_clk,      -- Connect to the 125MHz system clock
            reset      => sys_reset,    -- Connect to the system reset
            acl_data   => acl_data_int, -- Connect to the internal accelerometer data signal

            leds_out   => leds          -- Connect to the physical LED output pins
        );

    -- Note: The spi_busy_int signal is not directly used as an output
    -- in this top level, but it is used internally by the acl_led_indicator
    -- if you choose to modify it to show SPI busy status on an LED.
    -- Currently, acl_led_indicator uses acl_data != 0 to light LED0.

end architecture structural;
